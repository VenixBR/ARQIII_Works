module ControlPath (

);

endmodule 