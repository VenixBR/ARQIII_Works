module Top (

);

endmodule