module DataPath (

);

endmodule