module CLA (
    input  wire [15:0] A_i,
    input  wire [15:0] B_i,
    input  wire             Ci_i,
    output wire [15:0] S_o,
    output wire             Co_o
);

// Internal signals
wire g[0:15];
wire p[0:15];
wire c[0:15];
wire temp [0:15];

// Generate g and p functions
genvar i;
generate
    for(i=0 ; i<16 ; i=i+1)begin
        assign g[i] = A_i[i] & B_i[i];
        assign p[i] = A_i[i] ^ B_i[i];
    end
endgenerate

// Carries logic
assign c[0]  = Ci_i;
assign c[1]  = g[0]  | (p[0]  & c[0]);
assign c[2]  = g[1]  | (p[1]  & g[0])  | (p[1]  & p[0]  & c[0]) ;
assign c[3]  = g[2]  | (p[2]  & g[1])  | (p[2]  & p[1]  & g[0])  | (p[2]  & p[1]  & p[0]  & c[0]);
assign c[4]  = g[3]  | (p[3]  & g[2])  | (p[3]  & p[2]  & g[1])  | (p[3]  & p[2]  & p[1]  & g[0])  | (p[3]  & p[2]  & p[1]  & p[0]  & c[0]);
assign c[5]  = g[4]  | (p[4]  & g[3])  | (p[4]  & p[3]  & g[2])  | (p[4]  & p[3]  & p[2]  & g[1])  | (p[4]  & p[3]  & p[2]  & p[1]  & g[0])  | (p[4]  & p[3]  & p[2]  & p[1]  & p[0]  & c[0]);
assign c[6]  = g[5]  | (p[5]  & g[4])  | (p[5]  & p[4]  & g[3])  | (p[5]  & p[4]  & p[3]  & g[2])  | (p[5]  & p[4]  & p[3]  & p[2]  & g[1])  | (p[5]  & p[4]  & p[3]  & p[2]  & p[1]  & g[0]) | (p[5]  & p[4]  & p[3]  & p[2]  & p[1]  & p[0] & c[0]);
assign c[7]  = g[6]  | (p[6]  & g[5])  | (p[6]  & p[5]  & g[4])  | (p[6]  & p[5]  & p[4]  & g[3])  | (p[6]  & p[5]  & p[4]  & p[3]  & g[2])  | (p[6]  & p[5]  & p[4]  & p[3]  & p[2]  & g[1]) | (p[6]  & p[5]  & p[4]  & p[3]  & p[2]  & p[1] & g[0]) | (p[6]  & p[5]  & p[4]  & p[3]  & p[2]  & p[1] & p[0] & c[0]);
assign c[8]  = g[7]  | (p[7]  & g[6])  | (p[7]  & p[6]  & g[5])  | (p[7]  & p[6]  & p[5]  & g[4])  | (p[7]  & p[6]  & p[5]  & p[4]  & g[3])  | (p[7]  & p[6]  & p[5]  & p[4]  & p[3]  & g[2]) | (p[7]  & p[6]  & p[5]  & p[4]  & p[3]  & p[2] & g[1]) | (p[7]  & p[6]  & p[5]  & p[4]  & p[3]  & p[2] & p[1] & g[0]) | (p[7]  & p[6]  & p[5]  & p[4]  & p[3]  & p[2] & p[1] & p[0] & c[0]);
assign c[9]  = g[8]  | (p[8]  & g[7])  | (p[8]  & p[7]  & g[6])  | (p[8]  & p[7]  & p[6]  & g[5])  | (p[8]  & p[7]  & p[6]  & p[5]  & g[4])  | (p[8]  & p[7]  & p[6]  & p[5]  & p[4]  & g[3]) | (p[8]  & p[7]  & p[6]  & p[5]  & p[4]  & p[3] & g[2]) | (p[8]  & p[7]  & p[6]  & p[5]  & p[4]  & p[3] & p[2] & g[1]) | (p[8]  & p[7]  & p[6]  & p[5]  & p[4]  & p[3] & p[2] & p[1] & g[0]) | (p[8]  & p[7]  & p[6]  & p[5]  & p[4]  & p[3] & p[2] & p[1] & p[0] & c[0]);
assign c[10] = g[9]  | (p[9]  & g[8])  | (p[9]  & p[8]  & g[7])  | (p[9]  & p[8]  & p[7]  & g[6])  | (p[9]  & p[8]  & p[7]  & p[6]  & g[5])  | (p[9]  & p[8]  & p[7]  & p[6]  & p[5]  & g[4]) | (p[9]  & p[8]  & p[7]  & p[6]  & p[5]  & p[4] & g[3]) | (p[9]  & p[8]  & p[7]  & p[6]  & p[5]  & p[4] & p[3] & g[2]) | (p[9]  & p[8]  & p[7]  & p[6]  & p[5]  & p[4] & p[3] & p[2] & g[1]) | (p[9]  & p[8]  & p[7]  & p[6]  & p[5]  & p[4] & p[3] & p[2] & p[1] & g[0]) | (p[9]  & p[8]  & p[7]  & p[6]  & p[5]  & p[4] & p[3] & p[2] & p[1] & p[0] & c[0]);
assign c[11] = g[10] | (p[10] & g[9])  | (p[10] & p[9]  & g[8])  | (p[10] & p[9]  & p[8]  & g[7])  | (p[10] & p[9]  & p[8]  & p[7]  & g[6])  | (p[10] & p[9]  & p[8]  & p[7]  & p[6]  & g[5]) | (p[10] & p[9]  & p[8]  & p[7]  & p[6]  & p[5] & g[4]) | (p[10] & p[9]  & p[8]  & p[7]  & p[6]  & p[5] & p[4] & g[3]) | (p[10] & p[9]  & p[8]  & p[7]  & p[6]  & p[5] & p[4] & p[3] & g[2]) | (p[10] & p[9]  & p[8]  & p[7]  & p[6]  & p[5] & p[4] & p[3] & p[2] & g[1]) | (p[10] & p[9]  & p[8]  & p[7]  & p[6]  & p[5] & p[4] & p[3] & p[2] & p[1] & g[0]) | (p[10] & p[9]  & p[8]  & p[7]  & p[6]  & p[5] & p[4] & p[3] & p[2] & p[1] & p[0] & c[0]);
assign c[12] = g[11] | (p[11] & g[10]) | (p[11] & p[10] & g[9])  | (p[11] & p[10] & p[9]  & g[8])  | (p[11] & p[10] & p[9]  & p[8]  & g[7])  | (p[11] & p[10] & p[9]  & p[8]  & p[7]  & g[6]) | (p[11] & p[10] & p[9]  & p[8]  & p[7]  & p[6] & g[5]) | (p[11] & p[10] & p[9]  & p[8]  & p[7]  & p[6] & p[5] & g[4]) | (p[11] & p[10] & p[9]  & p[8]  & p[7]  & p[6] & p[5] & p[4] & g[3]) | (p[11] & p[10] & p[9]  & p[8]  & p[7]  & p[6] & p[5] & p[4] & p[3] & g[2]) | (p[11] & p[10] & p[9]  & p[8]  & p[7]  & p[6] & p[5] & p[4] & p[3] & p[2] & g[1]) | (p[11] & p[10] & p[9]  & p[8]  & p[7]  & p[6] & p[5] & p[4] & p[3] & p[2] & p[1] & g[0]) | (p[11] & p[10] & p[9]  & p[8]  & p[7]  & p[6] & p[5] & p[4] & p[3] & p[2] & p[1] & p[0] & c[0]);
assign c[13] = g[12] | (p[12] & g[11]) | (p[12] & p[11] & g[10]) | (p[12] & p[11] & p[10] & g[9])  | (p[12] & p[11] & p[10] & p[9]  & g[8])  | (p[12] & p[11] & p[10] & p[9]  & p[8]  & g[7]) | (p[12] & p[11] & p[10] & p[9]  & p[8]  & p[7] & g[6]) | (p[12] & p[11] & p[10] & p[9]  & p[8]  & p[7] & p[6] & g[5]) | (p[12] & p[11] & p[10] & p[9]  & p[8]  & p[7] & p[6] & p[5] & g[4]) | (p[12] & p[11] & p[10] & p[9]  & p[8]  & p[7] & p[6] & p[5] & p[4] & g[3]) | (p[12] & p[11] & p[10] & p[9]  & p[8]  & p[7] & p[6] & p[5] & p[4] & p[3] & g[2]) | (p[12] & p[11] & p[10] & p[9]  & p[8]  & p[7] & p[6] & p[5] & p[4] & p[3] & p[2] & g[1]) | (p[12] & p[11] & p[10] & p[9]  & p[8]  & p[7] & p[6] & p[5] & p[4] & p[3] & p[2] & p[1] & g[0]) | (p[12] & p[11] & p[10] & p[9]  & p[8]  & p[7] & p[6] & p[5] & p[4] & p[3] & p[2] & p[1] & p[0] & c[0]);
assign c[14] = g[13] | (p[13] & g[12]) | (p[13] & p[12] & g[11]) | (p[13] & p[12] & p[11] & g[10]) | (p[13] & p[12] & p[11] & p[10] & g[9])  | (p[13] & p[12] & p[11] & p[10] & p[9]  & g[8]) | (p[13] & p[12] & p[11] & p[10] & p[9]  & p[8] & g[7]) | (p[13] & p[12] & p[11] & p[10] & p[9]  & p[8] & p[7] & g[6]) | (p[13] & p[12] & p[11] & p[10] & p[9]  & p[8] & p[7] & p[6] & g[5]) | (p[13] & p[12] & p[11] & p[10] & p[9]  & p[8] & p[7] & p[6] & p[5] & g[4]) | (p[13] & p[12] & p[11] & p[10] & p[9]  & p[8] & p[7] & p[6] & p[5] & p[4] & g[3]) | (p[13] & p[12] & p[11] & p[10] & p[9]  & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & g[2]) | (p[13] & p[12] & p[11] & p[10] & p[9]  & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & p[2] & g[1]) | (p[13] & p[12] & p[11] & p[10] & p[9]  & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & p[2] & p[1] & g[0]) | (p[13] & p[12] & p[11] & p[10] & p[9]  & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & p[2] & p[1] & p[0] & c[0]);
assign c[15] = g[14] | (p[14] & g[13]) | (p[14] & p[13] & g[12]) | (p[14] & p[13] & p[12] & g[11]) | (p[14] & p[13] & p[12] & p[11] & g[10]) | (p[14] & p[13] & p[12] & p[11] & p[10] & g[9]) | (p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & g[8]) | (p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & g[7]) | (p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & g[6]) | (p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & g[5]) | (p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & g[4]) | (p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & g[3]) | (p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & g[2]) | (p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & p[2] & g[1]) | (p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & p[2] & p[1] & g[0]) | (p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & p[2] & p[1] & p[0] & c[0]);

assign Co_o = c[15];
// assign temp[0] = p[4] & p[3] & p[2];
// assign temp[1] = p[1] & p[0] & c[0];
// assign temp[3] = temp[1] & temp[2];
// assign temp[4] = g[4] | (p[4] & g[3]) | (p[4] & p[3] & g[2]) | (p[4] & p[3] & p[2] & g[1]) | (p[4] & p[3] & p[2] & p[1] & g[0]);
// assign c[5] = temp[4] | temp[3];

// Sums logic
assign S_o[0]  = p[0]  ^ c[0];
assign S_o[1]  = p[1]  ^ c[1];
assign S_o[2]  = p[2]  ^ c[2];
assign S_o[3]  = p[3]  ^ c[3];
assign S_o[4]  = p[4]  ^ c[4];
assign S_o[5]  = p[5]  ^ c[5];
assign S_o[6]  = p[6]  ^ c[6];
assign S_o[7]  = p[7]  ^ c[7];
assign S_o[8]  = p[8]  ^ c[8];
assign S_o[9]  = p[9]  ^ c[9];
assign S_o[10] = p[10] ^ c[10];
assign S_o[11] = p[11] ^ c[11];
assign S_o[12] = p[12] ^ c[12];
assign S_o[13] = p[13] ^ c[13];
assign S_o[14] = p[14] ^ c[14];
assign S_o[15] = p[15] ^ c[15];

endmodule